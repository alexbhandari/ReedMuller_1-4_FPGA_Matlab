module project (audio_in, aclk, clk, switch, audio_out);
	input [31:0] audio_in;
	input aclk;
	input clk;
	input [2:0] switch;
	output [31:0] audio_out;

	//quantize
	wire [9:0] audio_q = audio_in[31:22];
	
	//code blocks
	encode_corrupt_decode	ecd0	(	.audio_in(audio_q[9:5]),	.aclk(aclk), .clk(clk), .switch(switch), .audio_out(audio_out[31:27])	);
	encode_corrupt_decode	ecd1	(	.audio_in(audio_q[4:0]),	.aclk(aclk), .clk(clk), .switch(switch), .audio_out(audio_out[26:22])	);

	reg [0:15] e [0:696] = '{  16'b0000000000000000,
										16'b1000000000000000,
	                           16'b0100000000000000,
	                           16'b0010000000000000,
	                           16'b0001000000000000,
	                           16'b0000100000000000,
	                           16'b0000010000000000,
	                           16'b0000001000000000,
	                           16'b0000000100000000,
	                           16'b0000000010000000,
	                           16'b0000000001000000,
	                           16'b0000000000100000,
	                           16'b0000000000010000,
	                           16'b0000000000001000,
	                           16'b0000000000000100,
	                           16'b0000000000000010,
	                           16'b0000000000000001,
	                           16'b1100000000000000,
	                           16'b1010000000000000,
	                           16'b1001000000000000,
	                           16'b1000100000000000,
	                           16'b1000010000000000,
	                           16'b1000001000000000,
	                           16'b1000000100000000,
	                           16'b1000000010000000,
	                           16'b1000000001000000,
	                           16'b1000000000100000,
	                           16'b1000000000010000,
	                           16'b1000000000001000,
	                           16'b1000000000000100,
	                           16'b1000000000000010,
	                           16'b1000000000000001,
	                           16'b0110000000000000,
	                           16'b0101000000000000,
	                           16'b0100100000000000,
	                           16'b0100010000000000,
	                           16'b0100001000000000,
	                           16'b0100000100000000,
	                           16'b0100000010000000,
	                           16'b0100000001000000,
	                           16'b0100000000100000,
	                           16'b0100000000010000,
	                           16'b0100000000001000,
	                           16'b0100000000000100,
	                           16'b0100000000000010,
	                           16'b0100000000000001,
	                           16'b0011000000000000,
	                           16'b0010100000000000,
	                           16'b0010010000000000,
	                           16'b0010001000000000,
	                           16'b0010000100000000,
	                           16'b0010000010000000,
	                           16'b0010000001000000,
	                           16'b0010000000100000,
	                           16'b0010000000010000,
	                           16'b0010000000001000,
	                           16'b0010000000000100,
	                           16'b0010000000000010,
	                           16'b0010000000000001,
	                           16'b0001100000000000,
	                           16'b0001010000000000,
	                           16'b0001001000000000,
	                           16'b0001000100000000,
	                           16'b0001000010000000,
	                           16'b0001000001000000,
	                           16'b0001000000100000,
	                           16'b0001000000010000,
	                           16'b0001000000001000,
	                           16'b0001000000000100,
	                           16'b0001000000000010,
	                           16'b0001000000000001,
	                           16'b0000110000000000,
	                           16'b0000101000000000,
	                           16'b0000100100000000,
	                           16'b0000100010000000,
	                           16'b0000100001000000,
	                           16'b0000100000100000,
	                           16'b0000100000010000,
	                           16'b0000100000001000,
	                           16'b0000100000000100,
	                           16'b0000100000000010,
	                           16'b0000100000000001,
	                           16'b0000011000000000,
	                           16'b0000010100000000,
	                           16'b0000010010000000,
	                           16'b0000010001000000,
	                           16'b0000010000100000,
	                           16'b0000010000010000,
	                           16'b0000010000001000,
	                           16'b0000010000000100,
	                           16'b0000010000000010,
	                           16'b0000010000000001,
	                           16'b0000001100000000,
	                           16'b0000001010000000,
	                           16'b0000001001000000,
	                           16'b0000001000100000,
	                           16'b0000001000010000,
	                           16'b0000001000001000,
	                           16'b0000001000000100,
	                           16'b0000001000000010,
	                           16'b0000001000000001,
	                           16'b0000000110000000,
	                           16'b0000000101000000,
	                           16'b0000000100100000,
	                           16'b0000000100010000,
	                           16'b0000000100001000,
	                           16'b0000000100000100,
	                           16'b0000000100000010,
	                           16'b0000000100000001,
	                           16'b0000000011000000,
	                           16'b0000000010100000,
	                           16'b0000000010010000,
	                           16'b0000000010001000,
	                           16'b0000000010000100,
	                           16'b0000000010000010,
	                           16'b0000000010000001,
	                           16'b0000000001100000,
	                           16'b0000000001010000,
	                           16'b0000000001001000,
	                           16'b0000000001000100,
	                           16'b0000000001000010,
	                           16'b0000000001000001,
	                           16'b0000000000110000,
	                           16'b0000000000101000,
	                           16'b0000000000100100,
	                           16'b0000000000100010,
	                           16'b0000000000100001,
	                           16'b0000000000011000,
	                           16'b0000000000010100,
	                           16'b0000000000010010,
	                           16'b0000000000010001,
	                           16'b0000000000001100,
	                           16'b0000000000001010,
	                           16'b0000000000001001,
	                           16'b0000000000000110,
	                           16'b0000000000000101,
	                           16'b0000000000000011,
	                           16'b1110000000000000,
	                           16'b1101000000000000,
	                           16'b1100100000000000,
	                           16'b1100010000000000,
	                           16'b1100001000000000,
	                           16'b1100000100000000,
	                           16'b1100000010000000,
	                           16'b1100000001000000,
	                           16'b1100000000100000,
	                           16'b1100000000010000,
	                           16'b1100000000001000,
	                           16'b1100000000000100,
	                           16'b1100000000000010,
	                           16'b1100000000000001,
	                           16'b1011000000000000,
	                           16'b1010100000000000,
	                           16'b1010010000000000,
	                           16'b1010001000000000,
	                           16'b1010000100000000,
	                           16'b1010000010000000,
	                           16'b1010000001000000,
	                           16'b1010000000100000,
	                           16'b1010000000010000,
	                           16'b1010000000001000,
	                           16'b1010000000000100,
	                           16'b1010000000000010,
	                           16'b1010000000000001,
	                           16'b1001100000000000,
	                           16'b1001010000000000,
	                           16'b1001001000000000,
	                           16'b1001000100000000,
	                           16'b1001000010000000,
	                           16'b1001000001000000,
	                           16'b1001000000100000,
	                           16'b1001000000010000,
	                           16'b1001000000001000,
	                           16'b1001000000000100,
	                           16'b1001000000000010,
	                           16'b1001000000000001,
	                           16'b1000110000000000,
	                           16'b1000101000000000,
	                           16'b1000100100000000,
	                           16'b1000100010000000,
	                           16'b1000100001000000,
	                           16'b1000100000100000,
	                           16'b1000100000010000,
	                           16'b1000100000001000,
	                           16'b1000100000000100,
	                           16'b1000100000000010,
	                           16'b1000100000000001,
	                           16'b1000011000000000,
	                           16'b1000010100000000,
	                           16'b1000010010000000,
	                           16'b1000010001000000,
	                           16'b1000010000100000,
	                           16'b1000010000010000,
	                           16'b1000010000001000,
	                           16'b1000010000000100,
	                           16'b1000010000000010,
	                           16'b1000010000000001,
	                           16'b1000001100000000,
	                           16'b1000001010000000,
	                           16'b1000001001000000,
	                           16'b1000001000100000,
	                           16'b1000001000010000,
	                           16'b1000001000001000,
	                           16'b1000001000000100,
	                           16'b1000001000000010,
	                           16'b1000001000000001,
	                           16'b1000000110000000,
	                           16'b1000000101000000,
	                           16'b1000000100100000,
	                           16'b1000000100010000,
	                           16'b1000000100001000,
	                           16'b1000000100000100,
	                           16'b1000000100000010,
	                           16'b1000000100000001,
	                           16'b1000000011000000,
	                           16'b1000000010100000,
	                           16'b1000000010010000,
	                           16'b1000000010001000,
	                           16'b1000000010000100,
	                           16'b1000000010000010,
	                           16'b1000000010000001,
	                           16'b1000000001100000,
	                           16'b1000000001010000,
	                           16'b1000000001001000,
	                           16'b1000000001000100,
	                           16'b1000000001000010,
	                           16'b1000000001000001,
	                           16'b1000000000110000,
	                           16'b1000000000101000,
	                           16'b1000000000100100,
	                           16'b1000000000100010,
	                           16'b1000000000100001,
	                           16'b1000000000011000,
	                           16'b1000000000010100,
	                           16'b1000000000010010,
	                           16'b1000000000010001,
	                           16'b1000000000001100,
	                           16'b1000000000001010,
	                           16'b1000000000001001,
	                           16'b1000000000000110,
	                           16'b1000000000000101,
	                           16'b1000000000000011,
	                           16'b0111000000000000,
	                           16'b0110100000000000,
	                           16'b0110010000000000,
	                           16'b0110001000000000,
	                           16'b0110000100000000,
	                           16'b0110000010000000,
	                           16'b0110000001000000,
	                           16'b0110000000100000,
	                           16'b0110000000010000,
	                           16'b0110000000001000,
	                           16'b0110000000000100,
	                           16'b0110000000000010,
	                           16'b0110000000000001,
	                           16'b0101100000000000,
	                           16'b0101010000000000,
	                           16'b0101001000000000,
	                           16'b0101000100000000,
	                           16'b0101000010000000,
	                           16'b0101000001000000,
	                           16'b0101000000100000,
	                           16'b0101000000010000,
	                           16'b0101000000001000,
	                           16'b0101000000000100,
	                           16'b0101000000000010,
	                           16'b0101000000000001,
	                           16'b0100110000000000,
	                           16'b0100101000000000,
	                           16'b0100100100000000,
	                           16'b0100100010000000,
	                           16'b0100100001000000,
	                           16'b0100100000100000,
	                           16'b0100100000010000,
	                           16'b0100100000001000,
	                           16'b0100100000000100,
	                           16'b0100100000000010,
	                           16'b0100100000000001,
	                           16'b0100011000000000,
	                           16'b0100010100000000,
	                           16'b0100010010000000,
	                           16'b0100010001000000,
	                           16'b0100010000100000,
	                           16'b0100010000010000,
	                           16'b0100010000001000,
	                           16'b0100010000000100,
	                           16'b0100010000000010,
	                           16'b0100010000000001,
	                           16'b0100001100000000,
	                           16'b0100001010000000,
	                           16'b0100001001000000,
	                           16'b0100001000100000,
	                           16'b0100001000010000,
	                           16'b0100001000001000,
	                           16'b0100001000000100,
	                           16'b0100001000000010,
	                           16'b0100001000000001,
	                           16'b0100000110000000,
	                           16'b0100000101000000,
	                           16'b0100000100100000,
	                           16'b0100000100010000,
	                           16'b0100000100001000,
	                           16'b0100000100000100,
	                           16'b0100000100000010,
	                           16'b0100000100000001,
	                           16'b0100000011000000,
	                           16'b0100000010100000,
	                           16'b0100000010010000,
	                           16'b0100000010001000,
	                           16'b0100000010000100,
	                           16'b0100000010000010,
	                           16'b0100000010000001,
	                           16'b0100000001100000,
	                           16'b0100000001010000,
	                           16'b0100000001001000,
	                           16'b0100000001000100,
	                           16'b0100000001000010,
	                           16'b0100000001000001,
	                           16'b0100000000110000,
	                           16'b0100000000101000,
	                           16'b0100000000100100,
	                           16'b0100000000100010,
	                           16'b0100000000100001,
	                           16'b0100000000011000,
	                           16'b0100000000010100,
	                           16'b0100000000010010,
	                           16'b0100000000010001,
	                           16'b0100000000001100,
	                           16'b0100000000001010,
	                           16'b0100000000001001,
	                           16'b0100000000000110,
	                           16'b0100000000000101,
	                           16'b0100000000000011,
	                           16'b0011100000000000,
	                           16'b0011010000000000,
	                           16'b0011001000000000,
	                           16'b0011000100000000,
	                           16'b0011000010000000,
	                           16'b0011000001000000,
	                           16'b0011000000100000,
	                           16'b0011000000010000,
	                           16'b0011000000001000,
	                           16'b0011000000000100,
	                           16'b0011000000000010,
	                           16'b0011000000000001,
	                           16'b0010110000000000,
	                           16'b0010101000000000,
	                           16'b0010100100000000,
	                           16'b0010100010000000,
	                           16'b0010100001000000,
	                           16'b0010100000100000,
	                           16'b0010100000010000,
	                           16'b0010100000001000,
	                           16'b0010100000000100,
	                           16'b0010100000000010,
	                           16'b0010100000000001,
	                           16'b0010011000000000,
	                           16'b0010010100000000,
	                           16'b0010010010000000,
	                           16'b0010010001000000,
	                           16'b0010010000100000,
	                           16'b0010010000010000,
	                           16'b0010010000001000,
	                           16'b0010010000000100,
	                           16'b0010010000000010,
	                           16'b0010010000000001,
	                           16'b0010001100000000,
	                           16'b0010001010000000,
	                           16'b0010001001000000,
	                           16'b0010001000100000,
	                           16'b0010001000010000,
	                           16'b0010001000001000,
	                           16'b0010001000000100,
	                           16'b0010001000000010,
	                           16'b0010001000000001,
	                           16'b0010000110000000,
	                           16'b0010000101000000,
	                           16'b0010000100100000,
	                           16'b0010000100010000,
	                           16'b0010000100001000,
	                           16'b0010000100000100,
	                           16'b0010000100000010,
	                           16'b0010000100000001,
	                           16'b0010000011000000,
	                           16'b0010000010100000,
	                           16'b0010000010010000,
	                           16'b0010000010001000,
	                           16'b0010000010000100,
	                           16'b0010000010000010,
	                           16'b0010000010000001,
	                           16'b0010000001100000,
	                           16'b0010000001010000,
	                           16'b0010000001001000,
	                           16'b0010000001000100,
	                           16'b0010000001000010,
	                           16'b0010000001000001,
	                           16'b0010000000110000,
	                           16'b0010000000101000,
	                           16'b0010000000100100,
	                           16'b0010000000100010,
	                           16'b0010000000100001,
	                           16'b0010000000011000,
	                           16'b0010000000010100,
	                           16'b0010000000010010,
	                           16'b0010000000010001,
	                           16'b0010000000001100,
	                           16'b0010000000001010,
	                           16'b0010000000001001,
	                           16'b0010000000000110,
	                           16'b0010000000000101,
	                           16'b0010000000000011,
	                           16'b0001110000000000,
	                           16'b0001101000000000,
	                           16'b0001100100000000,
	                           16'b0001100010000000,
	                           16'b0001100001000000,
	                           16'b0001100000100000,
	                           16'b0001100000010000,
	                           16'b0001100000001000,
	                           16'b0001100000000100,
	                           16'b0001100000000010,
	                           16'b0001100000000001,
	                           16'b0001011000000000,
	                           16'b0001010100000000,
	                           16'b0001010010000000,
	                           16'b0001010001000000,
	                           16'b0001010000100000,
	                           16'b0001010000010000,
	                           16'b0001010000001000,
	                           16'b0001010000000100,
	                           16'b0001010000000010,
	                           16'b0001010000000001,
	                           16'b0001001100000000,
	                           16'b0001001010000000,
	                           16'b0001001001000000,
	                           16'b0001001000100000,
	                           16'b0001001000010000,
	                           16'b0001001000001000,
	                           16'b0001001000000100,
	                           16'b0001001000000010,
	                           16'b0001001000000001,
	                           16'b0001000110000000,
	                           16'b0001000101000000,
	                           16'b0001000100100000,
	                           16'b0001000100010000,
	                           16'b0001000100001000,
	                           16'b0001000100000100,
	                           16'b0001000100000010,
	                           16'b0001000100000001,
	                           16'b0001000011000000,
	                           16'b0001000010100000,
	                           16'b0001000010010000,
	                           16'b0001000010001000,
	                           16'b0001000010000100,
	                           16'b0001000010000010,
	                           16'b0001000010000001,
	                           16'b0001000001100000,
	                           16'b0001000001010000,
	                           16'b0001000001001000,
	                           16'b0001000001000100,
	                           16'b0001000001000010,
	                           16'b0001000001000001,
	                           16'b0001000000110000,
	                           16'b0001000000101000,
	                           16'b0001000000100100,
	                           16'b0001000000100010,
	                           16'b0001000000100001,
	                           16'b0001000000011000,
	                           16'b0001000000010100,
	                           16'b0001000000010010,
	                           16'b0001000000010001,
	                           16'b0001000000001100,
	                           16'b0001000000001010,
	                           16'b0001000000001001,
	                           16'b0001000000000110,
	                           16'b0001000000000101,
	                           16'b0001000000000011,
	                           16'b0000111000000000,
	                           16'b0000110100000000,
	                           16'b0000110010000000,
	                           16'b0000110001000000,
	                           16'b0000110000100000,
	                           16'b0000110000010000,
	                           16'b0000110000001000,
	                           16'b0000110000000100,
	                           16'b0000110000000010,
	                           16'b0000110000000001,
	                           16'b0000101100000000,
	                           16'b0000101010000000,
	                           16'b0000101001000000,
	                           16'b0000101000100000,
	                           16'b0000101000010000,
	                           16'b0000101000001000,
	                           16'b0000101000000100,
	                           16'b0000101000000010,
	                           16'b0000101000000001,
	                           16'b0000100110000000,
	                           16'b0000100101000000,
	                           16'b0000100100100000,
	                           16'b0000100100010000,
	                           16'b0000100100001000,
	                           16'b0000100100000100,
	                           16'b0000100100000010,
	                           16'b0000100100000001,
	                           16'b0000100011000000,
	                           16'b0000100010100000,
	                           16'b0000100010010000,
	                           16'b0000100010001000,
	                           16'b0000100010000100,
	                           16'b0000100010000010,
	                           16'b0000100010000001,
	                           16'b0000100001100000,
	                           16'b0000100001010000,
	                           16'b0000100001001000,
	                           16'b0000100001000100,
	                           16'b0000100001000010,
	                           16'b0000100001000001,
	                           16'b0000100000110000,
	                           16'b0000100000101000,
	                           16'b0000100000100100,
	                           16'b0000100000100010,
	                           16'b0000100000100001,
	                           16'b0000100000011000,
	                           16'b0000100000010100,
	                           16'b0000100000010010,
	                           16'b0000100000010001,
	                           16'b0000100000001100,
	                           16'b0000100000001010,
	                           16'b0000100000001001,
	                           16'b0000100000000110,
	                           16'b0000100000000101,
	                           16'b0000100000000011,
	                           16'b0000011100000000,
	                           16'b0000011010000000,
	                           16'b0000011001000000,
	                           16'b0000011000100000,
	                           16'b0000011000010000,
	                           16'b0000011000001000,
	                           16'b0000011000000100,
	                           16'b0000011000000010,
	                           16'b0000011000000001,
	                           16'b0000010110000000,
	                           16'b0000010101000000,
	                           16'b0000010100100000,
	                           16'b0000010100010000,
	                           16'b0000010100001000,
	                           16'b0000010100000100,
	                           16'b0000010100000010,
	                           16'b0000010100000001,
	                           16'b0000010011000000,
	                           16'b0000010010100000,
	                           16'b0000010010010000,
	                           16'b0000010010001000,
	                           16'b0000010010000100,
	                           16'b0000010010000010,
	                           16'b0000010010000001,
	                           16'b0000010001100000,
	                           16'b0000010001010000,
	                           16'b0000010001001000,
	                           16'b0000010001000100,
	                           16'b0000010001000010,
	                           16'b0000010001000001,
	                           16'b0000010000110000,
	                           16'b0000010000101000,
	                           16'b0000010000100100,
	                           16'b0000010000100010,
	                           16'b0000010000100001,
	                           16'b0000010000011000,
	                           16'b0000010000010100,
	                           16'b0000010000010010,
	                           16'b0000010000010001,
	                           16'b0000010000001100,
	                           16'b0000010000001010,
	                           16'b0000010000001001,
	                           16'b0000010000000110,
	                           16'b0000010000000101,
	                           16'b0000010000000011,
	                           16'b0000001110000000,
	                           16'b0000001101000000,
	                           16'b0000001100100000,
	                           16'b0000001100010000,
	                           16'b0000001100001000,
	                           16'b0000001100000100,
	                           16'b0000001100000010,
	                           16'b0000001100000001,
	                           16'b0000001011000000,
	                           16'b0000001010100000,
	                           16'b0000001010010000,
	                           16'b0000001010001000,
	                           16'b0000001010000100,
	                           16'b0000001010000010,
	                           16'b0000001010000001,
	                           16'b0000001001100000,
	                           16'b0000001001010000,
	                           16'b0000001001001000,
	                           16'b0000001001000100,
	                           16'b0000001001000010,
	                           16'b0000001001000001,
	                           16'b0000001000110000,
	                           16'b0000001000101000,
	                           16'b0000001000100100,
	                           16'b0000001000100010,
	                           16'b0000001000100001,
	                           16'b0000001000011000,
	                           16'b0000001000010100,
	                           16'b0000001000010010,
	                           16'b0000001000010001,
	                           16'b0000001000001100,
	                           16'b0000001000001010,
	                           16'b0000001000001001,
	                           16'b0000001000000110,
	                           16'b0000001000000101,
	                           16'b0000001000000011,
	                           16'b0000000111000000,
	                           16'b0000000110100000,
	                           16'b0000000110010000,
	                           16'b0000000110001000,
	                           16'b0000000110000100,
	                           16'b0000000110000010,
	                           16'b0000000110000001,
	                           16'b0000000101100000,
	                           16'b0000000101010000,
	                           16'b0000000101001000,
	                           16'b0000000101000100,
	                           16'b0000000101000010,
	                           16'b0000000101000001,
	                           16'b0000000100110000,
	                           16'b0000000100101000,
	                           16'b0000000100100100,
	                           16'b0000000100100010,
	                           16'b0000000100100001,
	                           16'b0000000100011000,
	                           16'b0000000100010100,
	                           16'b0000000100010010,
	                           16'b0000000100010001,
	                           16'b0000000100001100,
	                           16'b0000000100001010,
	                           16'b0000000100001001,
	                           16'b0000000100000110,
	                           16'b0000000100000101,
	                           16'b0000000100000011,
	                           16'b0000000011100000,
	                           16'b0000000011010000,
	                           16'b0000000011001000,
	                           16'b0000000011000100,
	                           16'b0000000011000010,
	                           16'b0000000011000001,
	                           16'b0000000010110000,
	                           16'b0000000010101000,
	                           16'b0000000010100100,
	                           16'b0000000010100010,
	                           16'b0000000010100001,
	                           16'b0000000010011000,
	                           16'b0000000010010100,
	                           16'b0000000010010010,
	                           16'b0000000010010001,
	                           16'b0000000010001100,
	                           16'b0000000010001010,
	                           16'b0000000010001001,
	                           16'b0000000010000110,
	                           16'b0000000010000101,
	                           16'b0000000010000011,
	                           16'b0000000001110000,
	                           16'b0000000001101000,
	                           16'b0000000001100100,
	                           16'b0000000001100010,
	                           16'b0000000001100001,
	                           16'b0000000001011000,
	                           16'b0000000001010100,
	                           16'b0000000001010010,
	                           16'b0000000001010001,
	                           16'b0000000001001100,
	                           16'b0000000001001010,
	                           16'b0000000001001001,
	                           16'b0000000001000110,
	                           16'b0000000001000101,
	                           16'b0000000001000011,
	                           16'b0000000000111000,
	                           16'b0000000000110100,
	                           16'b0000000000110010,
	                           16'b0000000000110001,
	                           16'b0000000000101100,
	                           16'b0000000000101010,
	                           16'b0000000000101001,
	                           16'b0000000000100110,
	                           16'b0000000000100101,
	                           16'b0000000000100011,
	                           16'b0000000000011100,
	                           16'b0000000000011010,
	                           16'b0000000000011001,
	                           16'b0000000000010110,
	                           16'b0000000000010101,
	                           16'b0000000000010011,
	                           16'b0000000000001110,
	                           16'b0000000000001101,
	                           16'b0000000000001011,
	                           16'b0000000000000111    };
										
   reg [0:15] eb [0:696] = '{ 11'b00000000000,
                              11'b11111100001,
                              11'b11100011101,
                              11'b10011011011,
                              11'b01010110111,
                              11'b00101101111,
                              11'b10000000000,
                              11'b01000000000,
                              11'b00100000000,
                              11'b00010000000,
                              11'b00001000000,
                              11'b00000100000,
                              11'b00000010000,
                              11'b00000001000,
                              11'b00000000100,
                              11'b00000000010,
                              11'b00000000001,
                              11'b00011111100,
                              11'b01100111010,
                              11'b10101010110,
                              11'b11010001110,
                              11'b01111100001,
                              11'b10111100001,
                              11'b11011100001,
                              11'b11101100001,
                              11'b11110100001,
                              11'b11111000001,
                              11'b11111110001,
                              11'b11111101001,
                              11'b11111100101,
                              11'b11111100011,
                              11'b11111100000,
                              11'b01111000110,
                              11'b10110101010,
                              11'b11001110010,
                              11'b01100011101,
                              11'b10100011101,
                              11'b11000011101,
                              11'b11110011101,
                              11'b11101011101,
                              11'b11100111101,
                              11'b11100001101,
                              11'b11100010101,
                              11'b11100011001,
                              11'b11100011111,
                              11'b11100011100,
                              11'b11001101100,
                              11'b10110110100,
                              11'b00011011011,
                              11'b11011011011,
                              11'b10111011011,
                              11'b10001011011,
                              11'b10010011011,
                              11'b10011111011,
                              11'b10011001011,
                              11'b10011010011,
                              11'b10011011111,
                              11'b10011011001,
                              11'b10011011010,
                              11'b01111011000,
                              11'b11010110111,
                              11'b00010110111,
                              11'b01110110111,
                              11'b01000110111,
                              11'b01011110111,
                              11'b01010010111,
                              11'b01010100111,
                              11'b01010111111,
                              11'b01010110011,
                              11'b01010110101,
                              11'b01010110110,
                              11'b10101101111,
                              11'b01101101111,
                              11'b00001101111,
                              11'b00111101111,
                              11'b00100101111,
                              11'b00101001111,
                              11'b00101111111,
                              11'b00101100111,
                              11'b00101101011,
                              11'b00101101101,
                              11'b00101101110,
                              11'b11000000000,
                              11'b10100000000,
                              11'b10010000000,
                              11'b10001000000,
                              11'b10000100000,
                              11'b10000010000,
                              11'b10000001000,
                              11'b10000000100,
                              11'b10000000010,
                              11'b10000000001,
                              11'b01100000000,
                              11'b01010000000,
                              11'b01001000000,
                              11'b01000100000,
                              11'b01000010000,
                              11'b01000001000,
                              11'b01000000100,
                              11'b01000000010,
                              11'b01000000001,
                              11'b00110000000,
                              11'b00101000000,
                              11'b00100100000,
                              11'b00100010000,
                              11'b00100001000,
                              11'b00100000100,
                              11'b00100000010,
                              11'b00100000001,
                              11'b00011000000,
                              11'b00010100000,
                              11'b00010010000,
                              11'b00010001000,
                              11'b00010000100,
                              11'b00010000010,
                              11'b00010000001,
                              11'b00001100000,
                              11'b00001010000,
                              11'b00001001000,
                              11'b00001000100,
                              11'b00001000010,
                              11'b00001000001,
                              11'b00000110000,
                              11'b00000101000,
                              11'b00000100100,
                              11'b00000100010,
                              11'b00000100001,
                              11'b00000011000,
                              11'b00000010100,
                              11'b00000010010,
                              11'b00000010001,
                              11'b00000001100,
                              11'b00000001010,
                              11'b00000001001,
                              11'b00000000110,
                              11'b00000000101,
                              11'b00000000011,
                              11'b10000100111,
                              11'b01001001011,
                              11'b00110010011,
                              11'b10011111100,
                              11'b01011111100,
                              11'b00111111100,
                              11'b00001111100,
                              11'b00010111100,
                              11'b00011011100,
                              11'b00011101100,
                              11'b00011110100,
                              11'b00011111000,
                              11'b00011111110,
                              11'b00011111101,
                              11'b00110001101,
                              11'b01001010101,
                              11'b11100111010,
                              11'b00100111010,
                              11'b01000111010,
                              11'b01110111010,
                              11'b01101111010,
                              11'b01100011010,
                              11'b01100101010,
                              11'b01100110010,
                              11'b01100111110,
                              11'b01100111000,
                              11'b01100111011,
                              11'b10000111001,
                              11'b00101010110,
                              11'b11101010110,
                              11'b10001010110,
                              11'b10111010110,
                              11'b10100010110,
                              11'b10101110110,
                              11'b10101000110,
                              11'b10101011110,
                              11'b10101010010,
                              11'b10101010100,
                              11'b10101010111,
                              11'b01010001110,
                              11'b10010001110,
                              11'b11110001110,
                              11'b11000001110,
                              11'b11011001110,
                              11'b11010101110,
                              11'b11010011110,
                              11'b11010000110,
                              11'b11010001010,
                              11'b11010001100,
                              11'b11010001111,
                              11'b00111100001,
                              11'b01011100001,
                              11'b01101100001,
                              11'b01110100001,
                              11'b01111000001,
                              11'b01111110001,
                              11'b01111101001,
                              11'b01111100101,
                              11'b01111100011,
                              11'b01111100000,
                              11'b10011100001,
                              11'b10101100001,
                              11'b10110100001,
                              11'b10111000001,
                              11'b10111110001,
                              11'b10111101001,
                              11'b10111100101,
                              11'b10111100011,
                              11'b10111100000,
                              11'b11001100001,
                              11'b11010100001,
                              11'b11011000001,
                              11'b11011110001,
                              11'b11011101001,
                              11'b11011100101,
                              11'b11011100011,
                              11'b11011100000,
                              11'b11100100001,
                              11'b11101000001,
                              11'b11101110001,
                              11'b11101101001,
                              11'b11101100101,
                              11'b11101100011,
                              11'b11101100000,
                              11'b11110000001,
                              11'b11110110001,
                              11'b11110101001,
                              11'b11110100101,
                              11'b11110100011,
                              11'b11110100000,
                              11'b11111010001,
                              11'b11111001001,
                              11'b11111000101,
                              11'b11111000011,
                              11'b11111000000,
                              11'b11111111001,
                              11'b11111110101,
                              11'b11111110011,
                              11'b11111110000,
                              11'b11111101101,
                              11'b11111101011,
                              11'b11111101000,
                              11'b11111100111,
                              11'b11111100100,
                              11'b11111100010,
                              11'b00101110001,
                              11'b01010101001,
                              11'b11111000110,
                              11'b00111000110,
                              11'b01011000110,
                              11'b01101000110,
                              11'b01110000110,
                              11'b01111100110,
                              11'b01111010110,
                              11'b01111001110,
                              11'b01111000010,
                              11'b01111000100,
                              11'b01111000111,
                              11'b10011000101,
                              11'b00110101010,
                              11'b11110101010,
                              11'b10010101010,
                              11'b10100101010,
                              11'b10111101010,
                              11'b10110001010,
                              11'b10110111010,
                              11'b10110100010,
                              11'b10110101110,
                              11'b10110101000,
                              11'b10110101011,
                              11'b01001110010,
                              11'b10001110010,
                              11'b11101110010,
                              11'b11011110010,
                              11'b11000110010,
                              11'b11001010010,
                              11'b11001100010,
                              11'b11001111010,
                              11'b11001110110,
                              11'b11001110000,
                              11'b11001110011,
                              11'b00100011101,
                              11'b01000011101,
                              11'b01110011101,
                              11'b01101011101,
                              11'b01100111101,
                              11'b01100001101,
                              11'b01100010101,
                              11'b01100011001,
                              11'b01100011111,
                              11'b01100011100,
                              11'b10000011101,
                              11'b10110011101,
                              11'b10101011101,
                              11'b10100111101,
                              11'b10100001101,
                              11'b10100010101,
                              11'b10100011001,
                              11'b10100011111,
                              11'b10100011100,
                              11'b11010011101,
                              11'b11001011101,
                              11'b11000111101,
                              11'b11000001101,
                              11'b11000010101,
                              11'b11000011001,
                              11'b11000011111,
                              11'b11000011100,
                              11'b11111011101,
                              11'b11110111101,
                              11'b11110001101,
                              11'b11110010101,
                              11'b11110011001,
                              11'b11110011111,
                              11'b11110011100,
                              11'b11101111101,
                              11'b11101001101,
                              11'b11101010101,
                              11'b11101011001,
                              11'b11101011111,
                              11'b11101011100,
                              11'b11100101101,
                              11'b11100110101,
                              11'b11100111001,
                              11'b11100111111,
                              11'b11100111100,
                              11'b11100000101,
                              11'b11100001001,
                              11'b11100001111,
                              11'b11100001100,
                              11'b11100010001,
                              11'b11100010111,
                              11'b11100010100,
                              11'b11100011011,
                              11'b11100011000,
                              11'b11100011110,
                              11'b11100000011,
                              11'b01001101100,
                              11'b10001101100,
                              11'b11101101100,
                              11'b11011101100,
                              11'b11000101100,
                              11'b11001001100,
                              11'b11001111100,
                              11'b11001100100,
                              11'b11001101000,
                              11'b11001101110,
                              11'b11001101101,
                              11'b00110110100,
                              11'b11110110100,
                              11'b10010110100,
                              11'b10100110100,
                              11'b10111110100,
                              11'b10110010100,
                              11'b10110100100,
                              11'b10110111100,
                              11'b10110110000,
                              11'b10110110110,
                              11'b10110110101,
                              11'b01011011011,
                              11'b00111011011,
                              11'b00001011011,
                              11'b00010011011,
                              11'b00011111011,
                              11'b00011001011,
                              11'b00011010011,
                              11'b00011011111,
                              11'b00011011001,
                              11'b00011011010,
                              11'b11111011011,
                              11'b11001011011,
                              11'b11010011011,
                              11'b11011111011,
                              11'b11011001011,
                              11'b11011010011,
                              11'b11011011111,
                              11'b11011011001,
                              11'b11011011010,
                              11'b10101011011,
                              11'b10110011011,
                              11'b10111111011,
                              11'b10111001011,
                              11'b10111010011,
                              11'b10111011111,
                              11'b10111011001,
                              11'b10111011010,
                              11'b10000011011,
                              11'b10001111011,
                              11'b10001001011,
                              11'b10001010011,
                              11'b10001011111,
                              11'b10001011001,
                              11'b10001011010,
                              11'b10010111011,
                              11'b10010001011,
                              11'b10010010011,
                              11'b10010011111,
                              11'b10010011001,
                              11'b10010011010,
                              11'b10011101011,
                              11'b10011110011,
                              11'b10011111111,
                              11'b10011111001,
                              11'b10011111010,
                              11'b10011000011,
                              11'b10011001111,
                              11'b10011001001,
                              11'b10011001010,
                              11'b10011010111,
                              11'b10011010001,
                              11'b10011010010,
                              11'b10011011101,
                              11'b10011011110,
                              11'b10011011000,
                              11'b11111011000,
                              11'b00111011000,
                              11'b01011011000,
                              11'b01101011000,
                              11'b01110011000,
                              11'b01111111000,
                              11'b01111001000,
                              11'b01111010000,
                              11'b01111011100,
                              11'b01111011010,
                              11'b01111011001,
                              11'b10010110111,
                              11'b11110110111,
                              11'b11000110111,
                              11'b11011110111,
                              11'b11010010111,
                              11'b11010100111,
                              11'b11010111111,
                              11'b11010110011,
                              11'b11010110101,
                              11'b11010110110,
                              11'b00110110111,
                              11'b00000110111,
                              11'b00011110111,
                              11'b00010010111,
                              11'b00010100111,
                              11'b00010111111,
                              11'b00010110011,
                              11'b00010110101,
                              11'b00010110110,
                              11'b01100110111,
                              11'b01111110111,
                              11'b01110010111,
                              11'b01110100111,
                              11'b01110111111,
                              11'b01110110011,
                              11'b01110110101,
                              11'b01110110110,
                              11'b01001110111,
                              11'b01000010111,
                              11'b01000100111,
                              11'b01000111111,
                              11'b01000110011,
                              11'b01000110101,
                              11'b01000110110,
                              11'b01011010111,
                              11'b01011100111,
                              11'b01011111111,
                              11'b01011110011,
                              11'b01011110101,
                              11'b01011110110,
                              11'b01010000111,
                              11'b01010011111,
                              11'b01010010011,
                              11'b01010010101,
                              11'b01010010110,
                              11'b01010101111,
                              11'b01010100011,
                              11'b01010100101,
                              11'b01010100110,
                              11'b01010111011,
                              11'b01010111101,
                              11'b01010111110,
                              11'b01010110001,
                              11'b01010110010,
                              11'b01010110100,
                              11'b11101101111,
                              11'b10001101111,
                              11'b10111101111,
                              11'b10100101111,
                              11'b10101001111,
                              11'b10101111111,
                              11'b10101100111,
                              11'b10101101011,
                              11'b10101101101,
                              11'b10101101110,
                              11'b01001101111,
                              11'b01111101111,
                              11'b01100101111,
                              11'b01101001111,
                              11'b01101111111,
                              11'b01101100111,
                              11'b01101101011,
                              11'b01101101101,
                              11'b01101101110,
                              11'b00011101111,
                              11'b00000101111,
                              11'b00001001111,
                              11'b00001111111,
                              11'b00001100111,
                              11'b00001101011,
                              11'b00001101101,
                              11'b00001101110,
                              11'b00110101111,
                              11'b00111001111,
                              11'b00111111111,
                              11'b00111100111,
                              11'b00111101011,
                              11'b00111101101,
                              11'b00111101110,
                              11'b00100001111,
                              11'b00100111111,
                              11'b00100100111,
                              11'b00100101011,
                              11'b00100101101,
                              11'b00100101110,
                              11'b00101011111,
                              11'b00101000111,
                              11'b00101001011,
                              11'b00101001101,
                              11'b00101001110,
                              11'b00101110111,
                              11'b00101111011,
                              11'b00101111101,
                              11'b00101111110,
                              11'b00101100011,
                              11'b00101100101,
                              11'b00101100110,
                              11'b00101101001,
                              11'b00101101010,
                              11'b00101101100,
                              11'b11100000000,
                              11'b11010000000,
                              11'b11001000000,
                              11'b11000100000,
                              11'b11000010000,
                              11'b11000001000,
                              11'b11000000100,
                              11'b11000000010,
                              11'b11000000001,
                              11'b10110000000,
                              11'b10101000000,
                              11'b10100100000,
                              11'b10100010000,
                              11'b10100001000,
                              11'b10100000100,
                              11'b10100000010,
                              11'b10100000001,
                              11'b10011000000,
                              11'b10010100000,
                              11'b10010010000,
                              11'b10010001000,
                              11'b10010000100,
                              11'b10010000010,
                              11'b10010000001,
                              11'b10001100000,
                              11'b10001010000,
                              11'b10001001000,
                              11'b10001000100,
                              11'b10001000010,
                              11'b10001000001,
                              11'b10000110000,
                              11'b10000101000,
                              11'b10000100100,
                              11'b10000100010,
                              11'b10000100001,
                              11'b10000011000,
                              11'b10000010100,
                              11'b10000010010,
                              11'b10000010001,
                              11'b10000001100,
                              11'b10000001010,
                              11'b10000001001,
                              11'b10000000110,
                              11'b10000000101,
                              11'b10000000011,
                              11'b01110000000,
                              11'b01101000000,
                              11'b01100100000,
                              11'b01100010000,
                              11'b01100001000,
                              11'b01100000100,
                              11'b01100000010,
                              11'b01100000001,
                              11'b01011000000,
                              11'b01010100000,
                              11'b01010010000,
                              11'b01010001000,
                              11'b01010000100,
                              11'b01010000010,
                              11'b01010000001,
                              11'b01001100000,
                              11'b01001010000,
                              11'b01001001000,
                              11'b01001000100,
                              11'b01001000010,
                              11'b01001000001,
                              11'b01000110000,
                              11'b01000101000,
                              11'b01000100100,
                              11'b01000100010,
                              11'b01000100001,
                              11'b01000011000,
                              11'b01000010100,
                              11'b01000010010,
                              11'b01000010001,
                              11'b01000001100,
                              11'b01000001010,
                              11'b01000001001,
                              11'b01000000110,
                              11'b01000000101,
                              11'b01000000011,
                              11'b00111000000,
                              11'b00110100000,
                              11'b00110010000,
                              11'b00110001000,
                              11'b00110000100,
                              11'b00110000010,
                              11'b00110000001,
                              11'b00101100000,
                              11'b00101010000,
                              11'b00101001000,
                              11'b00101000100,
                              11'b00101000010,
                              11'b00101000001,
                              11'b00100110000,
                              11'b00100101000,
                              11'b00100100100,
                              11'b00100100010,
                              11'b00100100001,
                              11'b00100011000,
                              11'b00100010100,
                              11'b00100010010,
                              11'b00100010001,
                              11'b00100001100,
                              11'b00100001010,
                              11'b00100001001,
                              11'b00100000110,
                              11'b00100000101,
                              11'b00100000011,
                              11'b00011100000,
                              11'b00011010000,
                              11'b00011001000,
                              11'b00011000100,
                              11'b00011000010,
                              11'b00011000001,
                              11'b00010110000,
                              11'b00010101000,
                              11'b00010100100,
                              11'b00010100010,
                              11'b00010100001,
                              11'b00010011000,
                              11'b00010010100,
                              11'b00010010010,
                              11'b00010010001,
                              11'b00010001100,
                              11'b00010001010,
                              11'b00010001001,
                              11'b00010000110,
                              11'b00010000101,
                              11'b00010000011,
                              11'b00001110000,
                              11'b00001101000,
                              11'b00001100100,
                              11'b00001100010,
                              11'b00001100001,
                              11'b00001011000,
                              11'b00001010100,
                              11'b00001010010,
                              11'b00001010001,
                              11'b00001001100,
                              11'b00001001010,
                              11'b00001001001,
                              11'b00001000110,
                              11'b00001000101,
                              11'b00001000011,
                              11'b00000111000,
                              11'b00000110100,
                              11'b00000110010,
                              11'b00000110001,
                              11'b00000101100,
                              11'b00000101010,
                              11'b00000101001,
                              11'b00000100110,
                              11'b00000100101,
                              11'b00000100011,
                              11'b00000011100,
                              11'b00000011010,
                              11'b00000011001,
                              11'b00000010110,
                              11'b00000010101,
                              11'b00000010011,
                              11'b00000001110,
                              11'b00000001101,
                              11'b00000001011,
                              11'b00000000111   };										

endmodule