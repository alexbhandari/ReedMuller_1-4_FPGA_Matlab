module project (audio_in, aclk, clk, audio_out);
	input [31:0] audio_in;
	input aclk;
	input clk;
	output [31:0] audio_out;

	//quantize
	wire [9:0] audio_q = audio_in[31:22];

	//generator is a 16x5 matrix
	reg [15:0] G [0:4] = '{		16'b1000011111100001,
										16'b0100011100011101,
										16'b0010010011011011,
										16'b0001001010110111,
										16'b0000100101101111 };

	//parity check is a 11x16 matrix
	reg [15:0] H [0:10] = '{	16'b1110010000000000,
										16'b1101001000000000,
										16'b1100100100000000,
										16'b1011000010000000,
										16'b1010100001000000,
										16'b1001100000100000,
										16'b0111000000010000,
										16'b0110100000001000,
										16'b0101100000000100,
										16'b0011100000000010,
										16'b1111100000000001	};

	reg [15:0] e [0:695] = '{  16'b1000000000000000,
	                           16'b0100000000000000,
	                           16'b0010000000000000,
	                           16'b0001000000000000,
	                           16'b0000100000000000,
	                           16'b0000010000000000,
	                           16'b0000001000000000,
	                           16'b0000000100000000,
	                           16'b0000000010000000,
	                           16'b0000000001000000,
	                           16'b0000000000100000,
	                           16'b0000000000010000,
	                           16'b0000000000001000,
	                           16'b0000000000000100,
	                           16'b0000000000000010,
	                           16'b0000000000000001,
	                           16'b1100000000000000,
	                           16'b1010000000000000,
	                           16'b1001000000000000,
	                           16'b1000100000000000,
	                           16'b1000010000000000,
	                           16'b1000001000000000,
	                           16'b1000000100000000,
	                           16'b1000000010000000,
	                           16'b1000000001000000,
	                           16'b1000000000100000,
	                           16'b1000000000010000,
	                           16'b1000000000001000,
	                           16'b1000000000000100,
	                           16'b1000000000000010,
	                           16'b1000000000000001,
	                           16'b0110000000000000,
	                           16'b0101000000000000,
	                           16'b0100100000000000,
	                           16'b0100010000000000,
	                           16'b0100001000000000,
	                           16'b0100000100000000,
	                           16'b0100000010000000,
	                           16'b0100000001000000,
	                           16'b0100000000100000,
	                           16'b0100000000010000,
	                           16'b0100000000001000,
	                           16'b0100000000000100,
	                           16'b0100000000000010,
	                           16'b0100000000000001,
	                           16'b0011000000000000,
	                           16'b0010100000000000,
	                           16'b0010010000000000,
	                           16'b0010001000000000,
	                           16'b0010000100000000,
	                           16'b0010000010000000,
	                           16'b0010000001000000,
	                           16'b0010000000100000,
	                           16'b0010000000010000,
	                           16'b0010000000001000,
	                           16'b0010000000000100,
	                           16'b0010000000000010,
	                           16'b0010000000000001,
	                           16'b0001100000000000,
	                           16'b0001010000000000,
	                           16'b0001001000000000,
	                           16'b0001000100000000,
	                           16'b0001000010000000,
	                           16'b0001000001000000,
	                           16'b0001000000100000,
	                           16'b0001000000010000,
	                           16'b0001000000001000,
	                           16'b0001000000000100,
	                           16'b0001000000000010,
	                           16'b0001000000000001,
	                           16'b0000110000000000,
	                           16'b0000101000000000,
	                           16'b0000100100000000,
	                           16'b0000100010000000,
	                           16'b0000100001000000,
	                           16'b0000100000100000,
	                           16'b0000100000010000,
	                           16'b0000100000001000,
	                           16'b0000100000000100,
	                           16'b0000100000000010,
	                           16'b0000100000000001,
	                           16'b0000011000000000,
	                           16'b0000010100000000,
	                           16'b0000010010000000,
	                           16'b0000010001000000,
	                           16'b0000010000100000,
	                           16'b0000010000010000,
	                           16'b0000010000001000,
	                           16'b0000010000000100,
	                           16'b0000010000000010,
	                           16'b0000010000000001,
	                           16'b0000001100000000,
	                           16'b0000001010000000,
	                           16'b0000001001000000,
	                           16'b0000001000100000,
	                           16'b0000001000010000,
	                           16'b0000001000001000,
	                           16'b0000001000000100,
	                           16'b0000001000000010,
	                           16'b0000001000000001,
	                           16'b0000000110000000,
	                           16'b0000000101000000,
	                           16'b0000000100100000,
	                           16'b0000000100010000,
	                           16'b0000000100001000,
	                           16'b0000000100000100,
	                           16'b0000000100000010,
	                           16'b0000000100000001,
	                           16'b0000000011000000,
	                           16'b0000000010100000,
	                           16'b0000000010010000,
	                           16'b0000000010001000,
	                           16'b0000000010000100,
	                           16'b0000000010000010,
	                           16'b0000000010000001,
	                           16'b0000000001100000,
	                           16'b0000000001010000,
	                           16'b0000000001001000,
	                           16'b0000000001000100,
	                           16'b0000000001000010,
	                           16'b0000000001000001,
	                           16'b0000000000110000,
	                           16'b0000000000101000,
	                           16'b0000000000100100,
	                           16'b0000000000100010,
	                           16'b0000000000100001,
	                           16'b0000000000011000,
	                           16'b0000000000010100,
	                           16'b0000000000010010,
	                           16'b0000000000010001,
	                           16'b0000000000001100,
	                           16'b0000000000001010,
	                           16'b0000000000001001,
	                           16'b0000000000000110,
	                           16'b0000000000000101,
	                           16'b0000000000000011,
	                           16'b1110000000000000,
	                           16'b1101000000000000,
	                           16'b1100100000000000,
	                           16'b1100010000000000,
	                           16'b1100001000000000,
	                           16'b1100000100000000,
	                           16'b1100000010000000,
	                           16'b1100000001000000,
	                           16'b1100000000100000,
	                           16'b1100000000010000,
	                           16'b1100000000001000,
	                           16'b1100000000000100,
	                           16'b1100000000000010,
	                           16'b1100000000000001,
	                           16'b1011000000000000,
	                           16'b1010100000000000,
	                           16'b1010010000000000,
	                           16'b1010001000000000,
	                           16'b1010000100000000,
	                           16'b1010000010000000,
	                           16'b1010000001000000,
	                           16'b1010000000100000,
	                           16'b1010000000010000,
	                           16'b1010000000001000,
	                           16'b1010000000000100,
	                           16'b1010000000000010,
	                           16'b1010000000000001,
	                           16'b1001100000000000,
	                           16'b1001010000000000,
	                           16'b1001001000000000,
	                           16'b1001000100000000,
	                           16'b1001000010000000,
	                           16'b1001000001000000,
	                           16'b1001000000100000,
	                           16'b1001000000010000,
	                           16'b1001000000001000,
	                           16'b1001000000000100,
	                           16'b1001000000000010,
	                           16'b1001000000000001,
	                           16'b1000110000000000,
	                           16'b1000101000000000,
	                           16'b1000100100000000,
	                           16'b1000100010000000,
	                           16'b1000100001000000,
	                           16'b1000100000100000,
	                           16'b1000100000010000,
	                           16'b1000100000001000,
	                           16'b1000100000000100,
	                           16'b1000100000000010,
	                           16'b1000100000000001,
	                           16'b1000011000000000,
	                           16'b1000010100000000,
	                           16'b1000010010000000,
	                           16'b1000010001000000,
	                           16'b1000010000100000,
	                           16'b1000010000010000,
	                           16'b1000010000001000,
	                           16'b1000010000000100,
	                           16'b1000010000000010,
	                           16'b1000010000000001,
	                           16'b1000001100000000,
	                           16'b1000001010000000,
	                           16'b1000001001000000,
	                           16'b1000001000100000,
	                           16'b1000001000010000,
	                           16'b1000001000001000,
	                           16'b1000001000000100,
	                           16'b1000001000000010,
	                           16'b1000001000000001,
	                           16'b1000000110000000,
	                           16'b1000000101000000,
	                           16'b1000000100100000,
	                           16'b1000000100010000,
	                           16'b1000000100001000,
	                           16'b1000000100000100,
	                           16'b1000000100000010,
	                           16'b1000000100000001,
	                           16'b1000000011000000,
	                           16'b1000000010100000,
	                           16'b1000000010010000,
	                           16'b1000000010001000,
	                           16'b1000000010000100,
	                           16'b1000000010000010,
	                           16'b1000000010000001,
	                           16'b1000000001100000,
	                           16'b1000000001010000,
	                           16'b1000000001001000,
	                           16'b1000000001000100,
	                           16'b1000000001000010,
	                           16'b1000000001000001,
	                           16'b1000000000110000,
	                           16'b1000000000101000,
	                           16'b1000000000100100,
	                           16'b1000000000100010,
	                           16'b1000000000100001,
	                           16'b1000000000011000,
	                           16'b1000000000010100,
	                           16'b1000000000010010,
	                           16'b1000000000010001,
	                           16'b1000000000001100,
	                           16'b1000000000001010,
	                           16'b1000000000001001,
	                           16'b1000000000000110,
	                           16'b1000000000000101,
	                           16'b1000000000000011,
	                           16'b0111000000000000,
	                           16'b0110100000000000,
	                           16'b0110010000000000,
	                           16'b0110001000000000,
	                           16'b0110000100000000,
	                           16'b0110000010000000,
	                           16'b0110000001000000,
	                           16'b0110000000100000,
	                           16'b0110000000010000,
	                           16'b0110000000001000,
	                           16'b0110000000000100,
	                           16'b0110000000000010,
	                           16'b0110000000000001,
	                           16'b0101100000000000,
	                           16'b0101010000000000,
	                           16'b0101001000000000,
	                           16'b0101000100000000,
	                           16'b0101000010000000,
	                           16'b0101000001000000,
	                           16'b0101000000100000,
	                           16'b0101000000010000,
	                           16'b0101000000001000,
	                           16'b0101000000000100,
	                           16'b0101000000000010,
	                           16'b0101000000000001,
	                           16'b0100110000000000,
	                           16'b0100101000000000,
	                           16'b0100100100000000,
	                           16'b0100100010000000,
	                           16'b0100100001000000,
	                           16'b0100100000100000,
	                           16'b0100100000010000,
	                           16'b0100100000001000,
	                           16'b0100100000000100,
	                           16'b0100100000000010,
	                           16'b0100100000000001,
	                           16'b0100011000000000,
	                           16'b0100010100000000,
	                           16'b0100010010000000,
	                           16'b0100010001000000,
	                           16'b0100010000100000,
	                           16'b0100010000010000,
	                           16'b0100010000001000,
	                           16'b0100010000000100,
	                           16'b0100010000000010,
	                           16'b0100010000000001,
	                           16'b0100001100000000,
	                           16'b0100001010000000,
	                           16'b0100001001000000,
	                           16'b0100001000100000,
	                           16'b0100001000010000,
	                           16'b0100001000001000,
	                           16'b0100001000000100,
	                           16'b0100001000000010,
	                           16'b0100001000000001,
	                           16'b0100000110000000,
	                           16'b0100000101000000,
	                           16'b0100000100100000,
	                           16'b0100000100010000,
	                           16'b0100000100001000,
	                           16'b0100000100000100,
	                           16'b0100000100000010,
	                           16'b0100000100000001,
	                           16'b0100000011000000,
	                           16'b0100000010100000,
	                           16'b0100000010010000,
	                           16'b0100000010001000,
	                           16'b0100000010000100,
	                           16'b0100000010000010,
	                           16'b0100000010000001,
	                           16'b0100000001100000,
	                           16'b0100000001010000,
	                           16'b0100000001001000,
	                           16'b0100000001000100,
	                           16'b0100000001000010,
	                           16'b0100000001000001,
	                           16'b0100000000110000,
	                           16'b0100000000101000,
	                           16'b0100000000100100,
	                           16'b0100000000100010,
	                           16'b0100000000100001,
	                           16'b0100000000011000,
	                           16'b0100000000010100,
	                           16'b0100000000010010,
	                           16'b0100000000010001,
	                           16'b0100000000001100,
	                           16'b0100000000001010,
	                           16'b0100000000001001,
	                           16'b0100000000000110,
	                           16'b0100000000000101,
	                           16'b0100000000000011,
	                           16'b0011100000000000,
	                           16'b0011010000000000,
	                           16'b0011001000000000,
	                           16'b0011000100000000,
	                           16'b0011000010000000,
	                           16'b0011000001000000,
	                           16'b0011000000100000,
	                           16'b0011000000010000,
	                           16'b0011000000001000,
	                           16'b0011000000000100,
	                           16'b0011000000000010,
	                           16'b0011000000000001,
	                           16'b0010110000000000,
	                           16'b0010101000000000,
	                           16'b0010100100000000,
	                           16'b0010100010000000,
	                           16'b0010100001000000,
	                           16'b0010100000100000,
	                           16'b0010100000010000,
	                           16'b0010100000001000,
	                           16'b0010100000000100,
	                           16'b0010100000000010,
	                           16'b0010100000000001,
	                           16'b0010011000000000,
	                           16'b0010010100000000,
	                           16'b0010010010000000,
	                           16'b0010010001000000,
	                           16'b0010010000100000,
	                           16'b0010010000010000,
	                           16'b0010010000001000,
	                           16'b0010010000000100,
	                           16'b0010010000000010,
	                           16'b0010010000000001,
	                           16'b0010001100000000,
	                           16'b0010001010000000,
	                           16'b0010001001000000,
	                           16'b0010001000100000,
	                           16'b0010001000010000,
	                           16'b0010001000001000,
	                           16'b0010001000000100,
	                           16'b0010001000000010,
	                           16'b0010001000000001,
	                           16'b0010000110000000,
	                           16'b0010000101000000,
	                           16'b0010000100100000,
	                           16'b0010000100010000,
	                           16'b0010000100001000,
	                           16'b0010000100000100,
	                           16'b0010000100000010,
	                           16'b0010000100000001,
	                           16'b0010000011000000,
	                           16'b0010000010100000,
	                           16'b0010000010010000,
	                           16'b0010000010001000,
	                           16'b0010000010000100,
	                           16'b0010000010000010,
	                           16'b0010000010000001,
	                           16'b0010000001100000,
	                           16'b0010000001010000,
	                           16'b0010000001001000,
	                           16'b0010000001000100,
	                           16'b0010000001000010,
	                           16'b0010000001000001,
	                           16'b0010000000110000,
	                           16'b0010000000101000,
	                           16'b0010000000100100,
	                           16'b0010000000100010,
	                           16'b0010000000100001,
	                           16'b0010000000011000,
	                           16'b0010000000010100,
	                           16'b0010000000010010,
	                           16'b0010000000010001,
	                           16'b0010000000001100,
	                           16'b0010000000001010,
	                           16'b0010000000001001,
	                           16'b0010000000000110,
	                           16'b0010000000000101,
	                           16'b0010000000000011,
	                           16'b0001110000000000,
	                           16'b0001101000000000,
	                           16'b0001100100000000,
	                           16'b0001100010000000,
	                           16'b0001100001000000,
	                           16'b0001100000100000,
	                           16'b0001100000010000,
	                           16'b0001100000001000,
	                           16'b0001100000000100,
	                           16'b0001100000000010,
	                           16'b0001100000000001,
	                           16'b0001011000000000,
	                           16'b0001010100000000,
	                           16'b0001010010000000,
	                           16'b0001010001000000,
	                           16'b0001010000100000,
	                           16'b0001010000010000,
	                           16'b0001010000001000,
	                           16'b0001010000000100,
	                           16'b0001010000000010,
	                           16'b0001010000000001,
	                           16'b0001001100000000,
	                           16'b0001001010000000,
	                           16'b0001001001000000,
	                           16'b0001001000100000,
	                           16'b0001001000010000,
	                           16'b0001001000001000,
	                           16'b0001001000000100,
	                           16'b0001001000000010,
	                           16'b0001001000000001,
	                           16'b0001000110000000,
	                           16'b0001000101000000,
	                           16'b0001000100100000,
	                           16'b0001000100010000,
	                           16'b0001000100001000,
	                           16'b0001000100000100,
	                           16'b0001000100000010,
	                           16'b0001000100000001,
	                           16'b0001000011000000,
	                           16'b0001000010100000,
	                           16'b0001000010010000,
	                           16'b0001000010001000,
	                           16'b0001000010000100,
	                           16'b0001000010000010,
	                           16'b0001000010000001,
	                           16'b0001000001100000,
	                           16'b0001000001010000,
	                           16'b0001000001001000,
	                           16'b0001000001000100,
	                           16'b0001000001000010,
	                           16'b0001000001000001,
	                           16'b0001000000110000,
	                           16'b0001000000101000,
	                           16'b0001000000100100,
	                           16'b0001000000100010,
	                           16'b0001000000100001,
	                           16'b0001000000011000,
	                           16'b0001000000010100,
	                           16'b0001000000010010,
	                           16'b0001000000010001,
	                           16'b0001000000001100,
	                           16'b0001000000001010,
	                           16'b0001000000001001,
	                           16'b0001000000000110,
	                           16'b0001000000000101,
	                           16'b0001000000000011,
	                           16'b0000111000000000,
	                           16'b0000110100000000,
	                           16'b0000110010000000,
	                           16'b0000110001000000,
	                           16'b0000110000100000,
	                           16'b0000110000010000,
	                           16'b0000110000001000,
	                           16'b0000110000000100,
	                           16'b0000110000000010,
	                           16'b0000110000000001,
	                           16'b0000101100000000,
	                           16'b0000101010000000,
	                           16'b0000101001000000,
	                           16'b0000101000100000,
	                           16'b0000101000010000,
	                           16'b0000101000001000,
	                           16'b0000101000000100,
	                           16'b0000101000000010,
	                           16'b0000101000000001,
	                           16'b0000100110000000,
	                           16'b0000100101000000,
	                           16'b0000100100100000,
	                           16'b0000100100010000,
	                           16'b0000100100001000,
	                           16'b0000100100000100,
	                           16'b0000100100000010,
	                           16'b0000100100000001,
	                           16'b0000100011000000,
	                           16'b0000100010100000,
	                           16'b0000100010010000,
	                           16'b0000100010001000,
	                           16'b0000100010000100,
	                           16'b0000100010000010,
	                           16'b0000100010000001,
	                           16'b0000100001100000,
	                           16'b0000100001010000,
	                           16'b0000100001001000,
	                           16'b0000100001000100,
	                           16'b0000100001000010,
	                           16'b0000100001000001,
	                           16'b0000100000110000,
	                           16'b0000100000101000,
	                           16'b0000100000100100,
	                           16'b0000100000100010,
	                           16'b0000100000100001,
	                           16'b0000100000011000,
	                           16'b0000100000010100,
	                           16'b0000100000010010,
	                           16'b0000100000010001,
	                           16'b0000100000001100,
	                           16'b0000100000001010,
	                           16'b0000100000001001,
	                           16'b0000100000000110,
	                           16'b0000100000000101,
	                           16'b0000100000000011,
	                           16'b0000011100000000,
	                           16'b0000011010000000,
	                           16'b0000011001000000,
	                           16'b0000011000100000,
	                           16'b0000011000010000,
	                           16'b0000011000001000,
	                           16'b0000011000000100,
	                           16'b0000011000000010,
	                           16'b0000011000000001,
	                           16'b0000010110000000,
	                           16'b0000010101000000,
	                           16'b0000010100100000,
	                           16'b0000010100010000,
	                           16'b0000010100001000,
	                           16'b0000010100000100,
	                           16'b0000010100000010,
	                           16'b0000010100000001,
	                           16'b0000010011000000,
	                           16'b0000010010100000,
	                           16'b0000010010010000,
	                           16'b0000010010001000,
	                           16'b0000010010000100,
	                           16'b0000010010000010,
	                           16'b0000010010000001,
	                           16'b0000010001100000,
	                           16'b0000010001010000,
	                           16'b0000010001001000,
	                           16'b0000010001000100,
	                           16'b0000010001000010,
	                           16'b0000010001000001,
	                           16'b0000010000110000,
	                           16'b0000010000101000,
	                           16'b0000010000100100,
	                           16'b0000010000100010,
	                           16'b0000010000100001,
	                           16'b0000010000011000,
	                           16'b0000010000010100,
	                           16'b0000010000010010,
	                           16'b0000010000010001,
	                           16'b0000010000001100,
	                           16'b0000010000001010,
	                           16'b0000010000001001,
	                           16'b0000010000000110,
	                           16'b0000010000000101,
	                           16'b0000010000000011,
	                           16'b0000001110000000,
	                           16'b0000001101000000,
	                           16'b0000001100100000,
	                           16'b0000001100010000,
	                           16'b0000001100001000,
	                           16'b0000001100000100,
	                           16'b0000001100000010,
	                           16'b0000001100000001,
	                           16'b0000001011000000,
	                           16'b0000001010100000,
	                           16'b0000001010010000,
	                           16'b0000001010001000,
	                           16'b0000001010000100,
	                           16'b0000001010000010,
	                           16'b0000001010000001,
	                           16'b0000001001100000,
	                           16'b0000001001010000,
	                           16'b0000001001001000,
	                           16'b0000001001000100,
	                           16'b0000001001000010,
	                           16'b0000001001000001,
	                           16'b0000001000110000,
	                           16'b0000001000101000,
	                           16'b0000001000100100,
	                           16'b0000001000100010,
	                           16'b0000001000100001,
	                           16'b0000001000011000,
	                           16'b0000001000010100,
	                           16'b0000001000010010,
	                           16'b0000001000010001,
	                           16'b0000001000001100,
	                           16'b0000001000001010,
	                           16'b0000001000001001,
	                           16'b0000001000000110,
	                           16'b0000001000000101,
	                           16'b0000001000000011,
	                           16'b0000000111000000,
	                           16'b0000000110100000,
	                           16'b0000000110010000,
	                           16'b0000000110001000,
	                           16'b0000000110000100,
	                           16'b0000000110000010,
	                           16'b0000000110000001,
	                           16'b0000000101100000,
	                           16'b0000000101010000,
	                           16'b0000000101001000,
	                           16'b0000000101000100,
	                           16'b0000000101000010,
	                           16'b0000000101000001,
	                           16'b0000000100110000,
	                           16'b0000000100101000,
	                           16'b0000000100100100,
	                           16'b0000000100100010,
	                           16'b0000000100100001,
	                           16'b0000000100011000,
	                           16'b0000000100010100,
	                           16'b0000000100010010,
	                           16'b0000000100010001,
	                           16'b0000000100001100,
	                           16'b0000000100001010,
	                           16'b0000000100001001,
	                           16'b0000000100000110,
	                           16'b0000000100000101,
	                           16'b0000000100000011,
	                           16'b0000000011100000,
	                           16'b0000000011010000,
	                           16'b0000000011001000,
	                           16'b0000000011000100,
	                           16'b0000000011000010,
	                           16'b0000000011000001,
	                           16'b0000000010110000,
	                           16'b0000000010101000,
	                           16'b0000000010100100,
	                           16'b0000000010100010,
	                           16'b0000000010100001,
	                           16'b0000000010011000,
	                           16'b0000000010010100,
	                           16'b0000000010010010,
	                           16'b0000000010010001,
	                           16'b0000000010001100,
	                           16'b0000000010001010,
	                           16'b0000000010001001,
	                           16'b0000000010000110,
	                           16'b0000000010000101,
	                           16'b0000000010000011,
	                           16'b0000000001110000,
	                           16'b0000000001101000,
	                           16'b0000000001100100,
	                           16'b0000000001100010,
	                           16'b0000000001100001,
	                           16'b0000000001011000,
	                           16'b0000000001010100,
	                           16'b0000000001010010,
	                           16'b0000000001010001,
	                           16'b0000000001001100,
	                           16'b0000000001001010,
	                           16'b0000000001001001,
	                           16'b0000000001000110,
	                           16'b0000000001000101,
	                           16'b0000000001000011,
	                           16'b0000000000111000,
	                           16'b0000000000110100,
	                           16'b0000000000110010,
	                           16'b0000000000110001,
	                           16'b0000000000101100,
	                           16'b0000000000101010,
	                           16'b0000000000101001,
	                           16'b0000000000100110,
	                           16'b0000000000100101,
	                           16'b0000000000100011,
	                           16'b0000000000011100,
	                           16'b0000000000011010,
	                           16'b0000000000011001,
	                           16'b0000000000010110,
	                           16'b0000000000010101,
	                           16'b0000000000010011,
	                           16'b0000000000001110,
	                           16'b0000000000001101,
	                           16'b0000000000001011,
	                           16'b0000000000000111    };

	encode_corrupt_decode	ecd0	(	.audio_in(audio_q[9:6]),	.aclk(aclk), .clk(clk), .audio_out(audio_out[31:27])	);
	encode_corrupt_decode	ecd1	(	.audio_in(audio_q[5:0]),	.aclk(aclk), .clk(clk), .audio_out(audio_out[26:22])	);

endmodule